/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_asiclab_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output reg  [7:0] uo_out,   // Dedicated outputs (changed to reg)
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    wire reset = ~rst_n;

    // Set unused IOs to 0
    assign uio_out = 8'b0;
    assign uio_oe  = 8'b0;

    // Prevent unused signal warnings
    wire _unused = &{ena, uio_in, clk, rst_n, 1'b0};

    // Sequential logic for uo_out
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            uo_out <= 8'b0;
        end else begin
            // Lower 4 bits: sum of ui_in[7:4] and ui_in[3:0]
            // Upper 4 bits: sum of ui_in and uio_in
            uo_out[3:0] <= ui_in[7:4] + ui_in[3:0];
            uo_out[7:4] <= (ui_in + uio_in)[7:4];
        end
    end

endmodule
